module ROM(
	input wire[15:0] address,
	output reg[5:0] data
);
	
	(* rom_style = "block" *)

	always @*
	case(address)
	16'h0000:data=6'b000000;
    16'h0001:data=6'b000000;
    16'h0002:data=6'b010100;
    16'h0003:data=6'b111000;
    16'h0004:data=6'b001010;
    16'h0005:data=6'b101000;
    16'h0006:data=6'b001001;
    16'h0007:data=6'b001011;
    16'h0008:data=6'b111001;
    16'h0009:data=6'b000100;
    16'h000a:data=6'b110000;
    16'h000b:data=6'b111010;
    16'h000c:data=6'b100010;
    16'h000d:data=6'b101011;
    16'h000e:data=6'b100100;
    16'h000f:data=6'b100010;
    16'h0010:data=6'b100011;
    16'h0011:data=6'b110001;
    16'h0012:data=6'b101000;
    16'h0013:data=6'b101010;
    16'h0014:data=6'b111000;
    16'h0015:data=6'b000011;
    16'h0016:data=6'b110110;
    16'h0017:data=6'b000001;
    16'h0018:data=6'b111000;
    16'h0019:data=6'b000011;
    16'h001a:data=6'b111000;
    16'h001b:data=6'b001010;
    16'h001c:data=6'b101000;
    16'h001d:data=6'b000011;
    16'h001e:data=6'b001000;
    16'h001f:data=6'b001000;
    16'h0020:data=6'b001001;
    16'h0021:data=6'b001011;
    16'h0022:data=6'b111001;
    16'h0023:data=6'b000100;
    16'h0024:data=6'b000100;
    16'h0025:data=6'b011000;
    16'h0026:data=6'b000011;
    16'h0027:data=6'b111000;
    16'h0028:data=6'b001010;
    16'h0029:data=6'b101000;
    16'h002a:data=6'b000101;
    16'h002b:data=6'b000000;
    16'h002c:data=6'b001000;
    16'h002d:data=6'b001001;
    16'h002e:data=6'b001011;
    16'h002f:data=6'b111001;
    16'h0030:data=6'b000100;
    16'h0031:data=6'b000101;
    16'h0032:data=6'b101000;
    16'h0033:data=6'b001000;
    16'h0034:data=6'b100010;
    16'h0035:data=6'b100011;
    16'h0036:data=6'b110001;
    16'h0037:data=6'b101000;
    16'h0038:data=6'b000110;
    16'h0039:data=6'b001011;
    16'h003a:data=6'b001000;
    16'h003b:data=6'b101010;
    16'h003c:data=6'b111000;
    16'h003d:data=6'b000011;
    16'h003e:data=6'b110110;
    16'h003f:data=6'b000111;
    16'h0040:data=6'b100000;
    16'h0041:data=6'b001001;
    16'h0042:data=6'b100100;
    16'h0043:data=6'b100010;
    16'h0044:data=6'b100011;
    16'h0045:data=6'b110001;
    16'h0046:data=6'b101000;
    16'h0047:data=6'b101010;
    16'h0048:data=6'b111000;
    16'h0049:data=6'b000011;
    16'h004a:data=6'b110110;
    16'h004b:data=6'b001000;
    16'h004c:data=6'b110000;
    16'h004d:data=6'b001011;
    16'h004e:data=6'b111000;
    16'h004f:data=6'b001010;
    16'h0050:data=6'b101000;
    16'h0051:data=6'b001001;
    16'h0052:data=6'b001011;
    16'h0053:data=6'b111001;
    16'h0054:data=6'b000100;
    16'h0055:data=6'b110000;
    16'h0056:data=6'b111010;
    16'h0057:data=6'b100010;
    16'h0058:data=6'b101011;
    16'h0059:data=6'b001010;
    16'h005a:data=6'b000000;
    16'h005b:data=6'b001001;
    16'h005c:data=6'b100100;
    16'h005d:data=6'b100010;
    16'h005e:data=6'b100011;
    16'h005f:data=6'b110001;
    16'h0060:data=6'b101000;
    16'h0061:data=6'b101010;
    16'h0062:data=6'b111000;
    16'h0063:data=6'b000011;
    16'h0064:data=6'b110110;
    16'h0065:data=6'b001011;
    16'h0066:data=6'b010000;
    16'h0067:data=6'b001011;
    16'h0068:data=6'b111000;
    16'h0069:data=6'b001010;
    16'h006a:data=6'b101000;
    16'h006b:data=6'b001001;
    16'h006c:data=6'b001011;
    16'h006d:data=6'b111001;
    16'h006e:data=6'b000100;
    16'h006f:data=6'b110000;
    16'h0070:data=6'b111010;
    16'h0071:data=6'b100010;
    16'h0072:data=6'b101011;
    16'h0073:data=6'b011001;
    16'h0074:data=6'b000000;
    16'h0075:data=6'b010100;
    16'h0076:data=6'b111000;
    16'h0077:data=6'b001010;
    16'h0078:data=6'b101000;
    16'h0079:data=6'b001001;
    16'h007a:data=6'b001011;
    16'h007b:data=6'b111001;
    16'h007c:data=6'b000100;
    16'h007d:data=6'b110000;
    16'h007e:data=6'b111010;
    16'h007f:data=6'b100010;
    16'h0080:data=6'b101011;
    16'h0081:data=6'b100100;
    16'h0082:data=6'b100010;
    16'h0083:data=6'b100011;
    16'h0084:data=6'b110001;
    16'h0085:data=6'b101000;
    16'h0086:data=6'b101010;
    16'h0087:data=6'b111000;
    16'h0088:data=6'b000011;
    16'h0089:data=6'b110110;
	default :data=6'b111111;
	endcase

	// reg[15:0] address_reg = 16'h0000;
	// assign address = address_reg;
	// initial begin
	// 	#10
	// 	$display("%b",data);
	// end
endmodule